
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity seniales is
    port(
        light_1 : in std_logic_vector(3 downto 0);
        light_2 : in std_logic_vector(3 downto 0);
        light_3 : in std_logic_vector(3 downto 0);
        led_no_1 : in std_logic;
        led_no_2 : in std_logic;
        led_no_3 : in std_logic;
        
        

    );
end seniales;